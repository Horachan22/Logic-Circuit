/*
===================================================================
Project Name    : デコーダ
File Name       : 2_1.v
Encoding        : UTF-8
Creation Date   : 2021/4/22
===================================================================
*/

module decoder(a, x);

	input [2:0]a;
	output [7:0]x;

	and(x[0], ~a[0], ~a[1], ~a[2]);
	and(x[1],  a[0], ~a[1], ~a[2]);
	and(x[2], ~a[0],  a[1], ~a[2]);
	and(x[3],  a[0],  a[1], ~a[2]);
	and(x[4], ~a[0], ~a[1],  a[2]);
	and(x[5],  a[0], ~a[1],  a[2]);
	and(x[6], ~a[0],  a[1],  a[2]);
	and(x[7],  a[0],  a[1],  a[2]);

endmodule
