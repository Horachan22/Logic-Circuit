/*
===================================================================
Project Name    : エンコーダ
File Name       : 2_2.v
Encoding        : UTF-8
Creation Date   : 2021/4/22
===================================================================
*/

module encoder(a, x);

	input [7:0]a;
	output [3:0]x;

	wire [6:0]P;

	// assign x[0] = ~a[0] & (a[1] | ~a[2] & ~a[1] & ~a[0] & (a[3] | ~a[4] & (a[5] | a[7] & a[6] & ~a[5])));
	assign x[0] = ~a[0] & (a[1] | ~a[2] & ~a[1] & ~a[0] & (a[3] | ~a[4] & (a[7] & a[6] | a[5])));
	assign x[1] = ~a[0] & ~a[1] & (a[2] | a[3] | ~a[4] & ~a[5] & (a[6] | a[7]));
	assign x[2] = ~(a[0] | a[1] | a[2] | a[3]) & (a[4] | a[5] | a[6] | a[7]);
	assign x[3] = a[0] | a[1] | a[2] | a[3] | a[4] | a[5] | a[6] | a[7];

endmodule
